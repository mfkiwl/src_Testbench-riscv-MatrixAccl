package datatypes;
import FixedPoint::*;

typedef FixedPoint#(10,6) DataType;
typedef UInt#(16) ImgWidth;
typedef FixedPoint#(10,6) CoeffType;
typedef UInt#(12) BramWidth;
typedef UInt#(6) BramLength;

endpackage
